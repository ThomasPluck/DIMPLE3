module circular_buffer #(
    parameter WIDTH=32,
    parameter SPINS=32
)

endmodule